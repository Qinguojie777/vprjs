module if(
    input   clk,
);
endmodule
